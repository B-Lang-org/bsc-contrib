package GenCMsg where

import GenCRepr
import Vector
import qualified List
import FIFOF
import Semi_FIFOF

ctobBFIFOSize :: Integer
ctobBFIFOSize = 128
btocBFIFOSize :: Integer
btocBFIFOSize = 2
ctobCFIFOSize :: Integer
ctobCFIFOSize = 16
btocCFIFOSize :: Integer
btocCFIFOSize = 128

class FIFOs fifos ctobBytes ctobCount btocBytes btocCount | fifos -> ctobBytes ctobCount btocBytes btocCount where
  mkFIFOs :: Vector ctobCount (Reg (UInt 8)) -> UInt 8 -> ByteList -> Action ->
             Vector btocCount (Reg (UInt 8)) -> (UInt 8 -> ByteList -> Action) ->
             Module (fifos, Rules)

  genCMsgTypeHeaderDcls :: fifos -> State (List String) String
  genCMsgTypeImplDcls :: fifos -> State (List String) String
  genCFIFOStructItems :: fifos -> String
  genCFIFOInitCredits :: fifos -> String
  genCFIFORestoreCredits :: fifos -> String
  genCFIFOCollectCredits :: fifos -> String
  genCFIFOEncode :: fifos -> Integer -> String
  genCFIFODecode :: fifos -> Integer -> String
  genCFIFOHeaderDcls :: fifos -> String -> String
  genCFIFOImplDcls :: fifos -> String -> String

instance (Generic a r, FIFOs' r bcb ncb bbc nbc) => FIFOs a bcb ncb bbc nbc where
  mkFIFOs ctobCredits ctobTag ctobBody deq btocCredits enq = do
    (fifos, rs) <- mkFIFOs' ctobCredits ctobTag ctobBody deq btocCredits enq
    return (to fifos, rs)

  genCMsgTypeHeaderDcls _ = genCMsgTypeHeaderDcls' (_ :: r)
  genCMsgTypeImplDcls _ = genCMsgTypeImplDcls' (_ :: r)
  genCFIFOStructItems _ = genCFIFOStructItems' (_ :: r)
  genCFIFOInitCredits _ = genCFIFOInitCredits' (_ :: r)
  genCFIFORestoreCredits _ = genCFIFORestoreCredits' (_ :: r)
  genCFIFOCollectCredits _ = genCFIFOCollectCredits' (_ :: r)
  genCFIFOEncode _ = genCFIFOEncode' (_ :: r)
  genCFIFODecode _ = genCFIFODecode' (_ :: r)
  genCFIFOHeaderDcls _ = genCFIFOHeaderDcls' (_ :: r)
  genCFIFOImplDcls _ = genCFIFOImplDcls' (_ :: r)

class FIFOs' fifos ctobBytes ctobCount btocBytes btocCount | fifos -> ctobBytes ctobCount btocBytes btocCount where
  mkFIFOs' :: Vector ctobCount (Reg (UInt 8)) -> UInt 8 -> ByteList -> Action ->
              Vector btocCount (Reg (UInt 8)) -> (UInt 8 -> ByteList -> Action) ->
              Module (fifos, Rules)

  genCMsgTypeHeaderDcls' :: fifos -> State (List String) String
  genCMsgTypeImplDcls' :: fifos -> State (List String) String
  genCFIFOStructItems' :: fifos -> String
  genCFIFOInitCredits' :: fifos -> String
  genCFIFORestoreCredits' :: fifos -> String
  genCFIFOCollectCredits' :: fifos -> String
  genCFIFOEncode' :: fifos -> Integer -> String
  genCFIFODecode' :: fifos -> Integer -> String
  genCFIFOHeaderDcls' :: fifos -> String -> String
  genCFIFOImplDcls' :: fifos -> String -> String

instance (FIFOs' a bcb ncb bbc nbc) => FIFOs' (Meta m a) bcb ncb bbc nbc where
  mkFIFOs' ctobCredits ctobTag ctobBody deq btocCredits enq = do
    (fifos, rs) <- mkFIFOs' ctobCredits ctobTag ctobBody deq btocCredits enq
    return (Meta fifos, rs)

  genCMsgTypeHeaderDcls' _ = genCMsgTypeHeaderDcls' (_ :: a)
  genCMsgTypeImplDcls' _ = genCMsgTypeImplDcls' (_ :: a)
  genCFIFOStructItems' _ = genCFIFOStructItems' (_ :: a)
  genCFIFOInitCredits' _ = genCFIFOInitCredits' (_ :: a)
  genCFIFORestoreCredits' _ = genCFIFORestoreCredits' (_ :: a)
  genCFIFOCollectCredits' _ = genCFIFOCollectCredits' (_ :: a)
  genCFIFOEncode' _ = genCFIFOEncode' (_ :: a)
  genCFIFODecode' _ = genCFIFODecode' (_ :: a)
  genCFIFOHeaderDcls' _ = genCFIFOHeaderDcls' (_ :: a)
  genCFIFOImplDcls' _ = genCFIFOImplDcls' (_ :: a)

instance (FIFOs' a bcb1 ncb1 bbc1 nbc1, FIFOs' b bcb2 ncb2 bbc2 nbc2,
          Max bcb1 bcb2 bcb, Max bbc1 bbc2 bbc,
          Add bcb1 pcb1 bcb, Add bcb2 pcb2 bcb, Add bbc1 pbc1 bbc, Add bbc2 pbc2 bbc, 
          Add ncb1 ncb2 ncb, Add nbc1 nbc2 nbc) =>
         FIFOs' (a, b) bcb ncb bbc nbc where
  mkFIFOs' ctobCredits ctobTag ctobBody deq btocCredits enq = do
    (fifos1, rs1) <- mkFIFOs'
      (take ctobCredits) ctobTag ctobBody deq 
      (take btocCredits) (\ btocTag btocBody -> enq btocTag btocBody)
    (fifos2, rs2) <- mkFIFOs'
      (takeTail ctobCredits) ctobTag ctobBody deq 
      (takeTail btocCredits) (\ btocTag btocBody -> enq btocTag btocBody)
    return ((fifos1, fifos2), rs1 <+ rs2)

  genCMsgTypeHeaderDcls' _ = liftM2 strConcat (genCMsgTypeHeaderDcls' (_ :: a)) (genCMsgTypeHeaderDcls' (_ :: b))
  genCMsgTypeImplDcls' _ = liftM2 strConcat (genCMsgTypeImplDcls' (_ :: a)) (genCMsgTypeImplDcls' (_ :: b))
  genCFIFOStructItems' _ = genCFIFOStructItems' (_ :: a) +++ genCFIFOStructItems' (_ :: b)
  genCFIFOInitCredits' _ = genCFIFOInitCredits' (_ :: a) +++ genCFIFOInitCredits' (_ :: b)
  genCFIFORestoreCredits' _ = genCFIFORestoreCredits' (_ :: a) +++ genCFIFORestoreCredits' (_ :: b)
  genCFIFOCollectCredits' _ = genCFIFOCollectCredits' (_ :: a) +++ genCFIFOCollectCredits' (_ :: b)
  genCFIFOEncode' _ nbc = genCFIFOEncode' (_ :: a) nbc +++ genCFIFOEncode' (_ :: b) nbc
  genCFIFODecode' _ ncb = genCFIFODecode' (_ :: a) ncb +++ genCFIFODecode' (_ :: b) ncb
  genCFIFOHeaderDcls' _ name = genCFIFOHeaderDcls' (_ :: a) name +++ genCFIFOHeaderDcls' (_ :: b) name
  genCFIFOImplDcls' _ name = genCFIFOImplDcls' (_ :: a) name +++ genCFIFOImplDcls' (_ :: b) name

instance FIFOs' () 0 0 0 0 where
  mkFIFOs' _ _ _ _ _ _ = return ((), emptyRules)

  genCMsgTypeHeaderDcls' _ = return ""
  genCMsgTypeImplDcls' _ = return ""
  genCFIFOStructItems' _ = ""
  genCFIFOInitCredits' _ = ""
  genCFIFORestoreCredits' _ = ""
  genCFIFOCollectCredits' _ = ""
  genCFIFOEncode' _ _ = ""
  genCFIFODecode' _ _ = ""
  genCFIFOHeaderDcls' _ _ = ""
  genCFIFOImplDcls' _ _ = ""

-- C to B
instance (GenCRepr a gcrBytes, GenAllCDecls a, Bits a bBits) =>
         FIFOs' (Meta (MetaField name i) (Conc (FIFOF_O a))) gcrBytes 1 0 0 where
  mkFIFOs' ctobCredits ctobTag ctobBody deq _ _ = do
    fifo :: FIFOF a
    fifo <- mkSizedFIFOF ctobBFIFOSize
    let credits :: Reg (UInt 8)
        credits = head ctobCredits

    let fifo_o = FIFOF_O {
      first = fifo.first;
      deq   = do { credits := credits + 1; fifo.deq };
      notEmpty = fifo.notEmpty;
    }

    let ruleName = "handle_ctob_" +++ stringOf name
    let rs =
          rules
            ruleName: when ctobTag == fromInteger (valueOf i) ==> do
              fifo.enq (unpackBytes ctobBody).fst
              deq
    
    return (Meta $ Conc fifo_o, rs)

  genCMsgTypeHeaderDcls' _ = genAllCHeaderDecls (_ :: a)
  genCMsgTypeImplDcls' _ = genAllCImplDecls (_ :: a)
  genCFIFOStructItems' _ =
    let (lType, rType) = genCType (_ :: a)
    in "\t" +++ lType +++ " " +++ stringOf name +++ "_buf[" +++ integerToString ctobCFIFOSize +++ "]" +++ rType +++ ";\n" +++
       "\tuint8_t " +++ stringOf name +++ "_head;\n" +++
       "\tuint8_t " +++ stringOf name +++ "_size;\n" +++
       "\tuint8_t " +++ stringOf name +++ "_credits;\n" +++
       "\n"
  genCFIFOInitCredits' _ = ""
  genCFIFORestoreCredits' _ =
    "\tstate->" +++ stringOf name +++ "_credits += buf[credits_index++];\n"
  genCFIFOCollectCredits' _ = ""
  genCFIFOEncode' _ btocCount =
    "\tif (state->" +++ stringOf name +++ "_size > 0 && state->" +++ stringOf name +++ "_credits > 0) {\n" +++
    "\t\tbuf[" +++ integerToString btocCount +++ "] = " +++ integerToString (valueOf i) +++ ";\n" +++
    "\t\tuint8_t head_index = state->" +++ stringOf name +++ "_head % " +++ integerToString ctobCFIFOSize +++ ";\n" +++
    "\t\tuint8_t *data_buf = buf + " +++ integerToString (btocCount + 1) +++ ", *pack_buf = data_buf;\n" +++
    "\t\t" +++ genCPack (_ :: a) ("state->" +++ stringOf name +++ "_buf[head_index]") "&pack_buf" +++ "\n" +++
    "\t\tstate->" +++ stringOf name +++ "_head++;\n" +++
    "\t\tstate->" +++ stringOf name +++ "_size--;\n" +++
    "\t\tstate->" +++ stringOf name +++ "_credits--;\n" +++
    "\t\treturn pack_buf - data_buf;\n" +++
    "\t}\n\n"
  genCFIFODecode' _ _ = ""

  genCFIFOHeaderDcls' _ ifaceName =
    let (lType, rType) = genCType (_ :: a)
    in "// Enqueue a " +++ stringOf name +++ " message to send.\n" +++
       "// Return 0 if failed (queue overflow) or 1 if success.\n" +++
       "_Bool enqueue_" +++ ifaceName +++ "_" +++ stringOf name +++ "(" +++ ifaceName +++ "_state *, " +++ lType +++ " " +++ rType +++ ");\n\n"

  genCFIFOImplDcls' _ ifaceName =
    let (lType, rType) = genCType (_ :: a)
    in "_Bool enqueue_" +++ ifaceName +++ "_" +++ stringOf name +++ "(" +++ ifaceName +++ "_state *state, " +++ lType +++ " msg" +++ rType +++ ") {\n" +++
       "\tif (state->" +++ stringOf name +++ "_size >= " +++ integerToString ctobCFIFOSize +++ ") return 0; \n" +++
       "\tuint8_t tail_index = (state->" +++ stringOf name +++ "_head + state->" +++ stringOf name +++ "_size) % " +++ integerToString ctobCFIFOSize +++ ";\n" +++
       "\tstate->" +++ stringOf name +++ "_buf[tail_index] = msg;\n" +++
       "\tstate->" +++ stringOf name +++ "_size++;\n" +++
       "\treturn 1;\n" +++
       "}\n\n"

-- B to C
instance (GenCRepr a gcrBytes, GenAllCDecls a, Bits a bBits) =>
         FIFOs' (Meta (MetaField name i) (Conc (FIFOF_I a))) 0 0 gcrBytes 1 where
  mkFIFOs' _ _ _ _ btocCredits enq = do
    fifo :: FIFOF a
    fifo <- mkSizedFIFOF btocBFIFOSize
    let credits :: Reg (UInt 8)
        credits = head btocCredits

    let ruleName = "handle_btoc_" +++ stringOf name
    let rs =
          rules
            ruleName: when True ==> do
              credits := credits - 1
              enq (fromInteger $ valueOf i) $ packBytes fifo.first
              fifo.deq

    return (Meta $ Conc $ to_FIFOF_I fifo, rs)

  genCMsgTypeHeaderDcls' _ = genAllCHeaderDecls (_ :: a)
  genCMsgTypeImplDcls' _ = genAllCImplDecls (_ :: a)
  genCFIFOStructItems' _ =
    let (lType, rType) = genCType (_ :: a)
    in "\t" +++ lType +++ " " +++ stringOf name +++ "_buf[" +++ integerToString btocCFIFOSize +++ "]" +++ rType +++ ";\n" +++
       "\tuint8_t " +++ stringOf name +++ "_head;\n" +++
       "\tuint8_t " +++ stringOf name +++ "_size;\n" +++
       "\tuint8_t " +++ stringOf name +++ "_credits;\n" +++
       "\n"
  genCFIFOInitCredits' _ =
    "\tstate->" +++ stringOf name +++ "_credits = " +++ integerToString btocCFIFOSize +++ ";\n"
  genCFIFORestoreCredits' _ = ""
  genCFIFOCollectCredits' _ =
    "\ttotal_credits += state->" +++ stringOf name +++ "_credits;\n" +++
    "\tbuf[credits_index++] = state->" +++ stringOf name +++ "_credits;\n" +++
    "\tstate->" +++ stringOf name +++ "_credits = 0;\n\n"
  genCFIFOEncode' _ _ = ""
  genCFIFODecode' _ ctobCount =
    "\tif (buf[" +++ integerToString ctobCount +++ "] == " +++ integerToString (valueOf i) +++ ") {\n" +++
    "\t\tuint8_t tail_index = (state->" +++ stringOf name +++ "_head + state->" +++ stringOf name +++ "_size) % " +++ integerToString ctobCFIFOSize +++ ";\n" +++
    "\t\tuint8_t *data_buf = buf + " +++ integerToString (ctobCount + 1) +++ ";\n" +++
    "\t\t" +++ genCUnpack (_ :: a) ("state->" +++ stringOf name +++ "_buf[tail_index]") "&data_buf" +++ "\n" +++
    "\t\tstate->" +++ stringOf name +++ "_size++;\n" +++
    "\t\treturn 1;\n" +++
    "\t}\n\n"
  genCFIFODecode' _ _ = ""

  genCFIFOHeaderDcls' _ ifaceName =
    let (lType, rType) = genCType (_ :: a)
    in "// Dequeue a recieved " +++ stringOf name +++ " message.\n" +++
       "// Return 0 if failed (none available) or 1 if success.\n" +++
       "_Bool dequeue_" +++ ifaceName +++ "_" +++ stringOf name +++ "(" +++ ifaceName +++ "_state *, " +++ lType +++ " *" +++ rType +++ ");\n\n"

  genCFIFOImplDcls' _ ifaceName =
    let (lType, rType) = genCType (_ :: a)
    in "_Bool dequeue_" +++ ifaceName +++ "_" +++ stringOf name +++ "(" +++ ifaceName +++ "_state *state, " +++ lType +++ " *msg" +++ rType +++ ") {\n" +++
       "\tif (state->" +++ stringOf name +++ "_size == 0) return 0; \n" +++
       "\tuint8_t head_index = state->" +++ stringOf name +++ "_head % " +++ integerToString ctobCFIFOSize +++ ";\n" +++
       "\t*msg = state->" +++ stringOf name +++ "_buf[head_index];\n" +++
       "\tstate->" +++ stringOf name +++ "_head++;\n" +++
       "\tstate->" +++ stringOf name +++ "_size--;\n" +++
       "\tstate->" +++ stringOf name +++ "_credits++;\n" +++
       "\treturn 1;\n" +++
       "}\n\n"

interface MsgManager fifos ctobBytes btocBytes =
  fifos :: fifos
  putCToB :: Vector ctobBytes (Bit 8) -> Action
  getBToC :: ActionValue (UInt (TLog (TAdd 1 btocBytes)), Vector btocBytes (Bit 8))

class GenCMsg fifos ctobBytes btocBytes | fifos -> ctobBytes btocBytes where
  mkMsgManager :: Module (MsgManager fifos ctobBytes btocBytes)
  genCMsgHeaderDecls :: fifos -> State (List String) String
  genCMsgImplDecls :: fifos -> State (List String) String

instance (FIFOs fifos ctobBytes ctobCount btocBytes btocCount,
          Add btocCount 1 ctobHead, Add ctobHead ctobBytes ctobTotalBytes,
          Add btocCount ctobRest ctobTotalBytes,
          Add ctobCount 1 btocHead, Add btocHead btocBytes btocTotalBytes,
          Generic fifos (Meta (MetaData name pkg ta 1) r)) =>
         GenCMsg fifos ctobTotalBytes btocTotalBytes where
  mkMsgManager = module
    ctobMsgs :: FIFOF (Vector ctobTotalBytes (Bit 8))
    ctobMsgs <- mkFIFOF

    ctobCredits :: Vector ctobCount (Reg (UInt 8))
    ctobCredits <- replicateM $ mkReg $ fromInteger ctobBFIFOSize

    btocMsgs :: FIFOF (UInt (TLog (TAdd 1 btocTotalBytes)), Vector btocTotalBytes (Bit 8))
    btocMsgs <- mkFIFOF

    btocCredits :: Vector btocCount (Reg (UInt 8))
    btocCredits <- replicateM $ mkReg 0

    let ctobTag :: UInt 8
        ctobTag = unpack $ head ((drop ctobMsgs.first) :: Vector ctobHead (Bit 8))
    let ctobBody :: ByteList
        ctobBody = toList ((takeTail ctobMsgs.first) :: Vector ctobBytes (Bit 8))
    let deq :: Action
        deq = do
          zipWithM_ (\ cr c -> writeReg cr (cr + Prelude.unpack c)) btocCredits (take ctobMsgs.first)
          ctobMsgs.deq
    let enq :: UInt 8 -> ByteList -> Action
        enq btocTag btocBody = do
          mapM_ (flip writeReg 0) ctobCredits
          let packedCredits :: (Vector ctobCount (Bit 8))
              packedCredits = map (\ c -> Prelude.pack (c :: Reg (UInt 8))) ctobCredits
          let packedBody :: (Vector btocBytes (Bit 8))
              packedBody = toVector
                (btocBody `List.append` List.replicate (valueOf btocBytes - List.length btocBody) 0)
          btocMsgs.enq
            (fromInteger $ valueOf btocHead + List.length btocBody,
             packedCredits `append` (Prelude.pack btocTag :> packedBody))
    (fifos, rs) :: (fifos, Rules) <-
        mkFIFOs ctobCredits ctobTag ctobBody deq btocCredits enq

    let creditsOnlyTag = fromInteger $ valueOf ctobCount + valueOf btocCount
    let handleCreditsOnly =
          rules
             "handle_ctob_credits_only": when any (\ c -> readReg c > 0) ctobCredits ==> enq creditsOnlyTag List.nil
             "handle_btoc_credits_only": when ctobTag == creditsOnlyTag ==> deq
    addRules $ rs <+ handleCreditsOnly

    interface
      fifos = fifos
      putCToB = ctobMsgs.enq
      getBToC = do btocMsgs.deq; return btocMsgs.first

  genCMsgHeaderDecls _ = do
    deps <- genCMsgTypeHeaderDcls (_ :: fifos)
    let structItems = genCFIFOStructItems (_ :: fifos)
    return $ deps +++
      "typedef struct " +++ stringOf name +++ "_state {\n" +++
      structItems +++
      "} " +++ stringOf name +++ "_state;\n" +++
      "enum {\n" +++
      "\tsize_ctob_" +++ stringOf name +++ " = " +++ integerToString (valueOf ctobTotalBytes) +++ ",\n" +++
      "\tsize_btoc_" +++ stringOf name +++ " = " +++ integerToString (valueOf btocTotalBytes) +++ ",\n" +++
      "};\n\n" +++
      "// Initialize a message state struct.\n" +++
      "void init_" +++ stringOf name +++ "(" +++ stringOf name +++ "_state *);\n\n" +++
      "// Select and pack an available message.\n" +++
      "// Returns the size of the encoded message, or 0 if there is no message to send.\n" +++
      "size_t encode_" +++ stringOf name +++ "(" +++ stringOf name +++ "_state *, uint8_t buf[size_ctob_" +++ stringOf name +++ "]);\n\n" +++
      "// Unpack an incoming message.\n" +++
      "// Returns 1 if the message had a payload, or 0 if it is credits-only.\n" +++
      "_Bool decode_" +++ stringOf name +++ "(" +++ stringOf name +++ "_state *, uint8_t buf[size_btoc_" +++ stringOf name +++ "]);\n\n" +++
      genCFIFOHeaderDcls (_ :: fifos) (stringOf name) +++
      "\n"

  genCMsgImplDecls _ = do
    deps <- genCMsgTypeImplDcls (_ :: fifos)
    return $ deps +++
      "void init_" +++ stringOf name +++ "(" +++ stringOf name +++ "_state *state) {\n" +++
      "\tmemset(state, 0, sizeof(" +++ stringOf name +++ "_state));\n" +++
      genCFIFOInitCredits (_ :: fifos) +++
      "}\n\n" +++
      "size_t encode_" +++ stringOf name +++ "(" +++ stringOf name +++ "_state *state , uint8_t buf[size_ctob_" +++ stringOf name +++ "]) {\n" +++
      "\tuint32_t credits_index = 0;\n" +++
      "\tuint32_t total_credits = 0;\n" +++
      "\t\n" +++
      genCFIFOCollectCredits (_ :: fifos) +++
      genCFIFOEncode (_ :: fifos) (valueOf btocCount) +++
      "\t\n" +++
      "\tif (total_credits > 0) {\n" +++
      "\t\tbuf[" +++ integerToString (valueOf btocCount) +++ "] = " +++ integerToString (valueOf btocCount + valueOf ctobCount) +++ ";\n" +++
      "\t\treturn " +++ integerToString (valueOf btocCount + 1) +++ ";\n" +++
      "\t}\n" +++
      "\t\n" +++
      "\treturn 0; // Nothing to send\n" +++
      "}\n\n" +++
      "_Bool decode_" +++ stringOf name +++ "(" +++ stringOf name +++ "_state *state , uint8_t buf[size_btoc_" +++ stringOf name +++ "]) {\n" +++
      "\tuint32_t credits_index = 0;\n" +++
      genCFIFORestoreCredits (_ :: fifos) +++
      "\t\n" +++
      genCFIFODecode (_ :: fifos) (valueOf ctobCount) +++
      "\t\n" +++
      "\treturn 0; // Message is credits-only\n" +++
      "}\n\n" +++
      genCFIFOImplDcls (_ :: fifos) (stringOf name) +++
      "\n"

-- Driver to all write C declarations for a fifo interface
writeCMsgDecls :: (GenCMsg fifos ctobBytes btocBytes) => String -> fifos -> Module Empty
writeCMsgDecls baseName proxy = do
  let headerName = (baseName +++ ".h")
  let implName = (baseName +++ ".c")
  let headerContents =
        "#include <stdint.h>\n\n\n" +++
        (runState (genCMsgHeaderDecls proxy) List.nil).fst
  let implContents =
        "#include <stdlib.h>\n#include <string.h>\n\n#include \"" +++ headerName +++ "\"\n\n\n" +++
        (runState (genCMsgImplDecls proxy) List.nil).fst
  stdout <- openFile "/dev/stdout" WriteMode
  h <- openFile headerName WriteMode
  hPutStr h headerContents
  hClose h
  hPutStrLn stdout ("Message library header file created: " +++ headerName)
  c <- openFile implName WriteMode
  hPutStr c implContents
  hClose c
  hPutStrLn stdout ("Message library C implementation file created: " +++ implName)
  hClose stdout
