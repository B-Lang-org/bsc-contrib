////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause
//
////////////////////////////////////////////////////////////////////////////////
//  Filename      : XilinxUtils.bsv
//  Description   : Xilinx evaluation board utilities
////////////////////////////////////////////////////////////////////////////////
package XilinxUtils;

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import DIPSwitch        ::*;
import ButtonController ::*;
import LEDController    ::*;
import LCDController    ::*;
import DVIController    ::*;
import GPIOController   ::*;
import HDMIController   ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export DIPSwitch        ::*;
export ButtonController ::*;
export LEDController    ::*;
export LCDController    ::*;
export DVIController    ::*;
export GPIOController   ::*;
export HDMIController   ::*;

endpackage: XilinxUtils
