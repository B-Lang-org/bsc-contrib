
import "BDPI" function Bit#(48) getInstr(UInt#(8) ic);
import "BDPI" function Bit#(8) putResult(Bit#(48) res);

