// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause

package FPGA_Misc;

// Imports
import ClkCtrlServer     ::*;
import DDR3              ::*;
import DDR4              ::*;
import I2C               ::*;
import PCIE              ::*;
import PTMClocks         ::*;
import RS232             ::*;
import Video             ::*;

// Exports
export ClkCtrlServer     ::*;
export DDR3              ::*;
export DDR4              ::*;
export I2C               ::*;
export PCIE              ::*;
export PTMClocks         ::*;
export RS232             ::*;
export Video             ::*;

endpackage: FPGA_Misc
