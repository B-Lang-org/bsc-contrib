package Test where

import GenCRepr
import TestFn
import CShow

struct Foo =
  x :: UInt 8
  y :: Int 16
  z :: Bit 256

struct Bar =
  b :: Bool
  bs :: Bit 13
  f :: Foo

struct Baz = {}

data Qux = QA (UInt 16) | QB (UInt 8) | QC (UInt 32) --QF Foo | QFB Foo Bar | Q | QI { x :: Int 8; y :: Int 8} | QU { u :: UInt 16 }

struct Thing =
  x :: UInt 8
  y :: UInt 8
  z :: Int 16

struct ThingMsg =
  thing :: Thing
  swapXY :: Bool
  deltaZ :: Int 8

actTestThing :: ThingMsg -> Action
actTestThing tm = do
  $display (cshow tm)
  let input = GenCRepr.pack tm
  $display (cshow input)
  let output = toByteList $ test_fn $ fromByteList input
  $display (cshow output)
  let (res, _) = (GenCRepr.unpack output) :: (Thing, ByteList)
  $display (cshow res)

{-# verilog mkTest #-}
mkTest :: Module Empty
mkTest = module
  -- writeCDecls "test" ((error "proxy") :: (Foo, Bar, Baz, Qux, Thing, ThingMsg))
  writeCDecls "test" ((error "proxy") :: Qux)

  rules
    when True ==> do
      actTestThing (ThingMsg {thing=Thing {x=1; y=2; z=1234;}; swapXY=False; deltaZ=8;})
      actTestThing (ThingMsg {thing=Thing {x=1; y=2; z=1234;}; swapXY=True; deltaZ=negate 8;})
      $finish
