// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause

package TLM3;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import TLM3Api::*;
import TLM3BRAM::*;
import TLM3CBusAdapter::*;
import TLM3Defines::*;
import TLM3Limit::*;
import TLM3Reorder::*;
import TLM3FlowControl::*;
import TLM3Ram::*;
import TLM3ReadWriteRam::*;
import TLM3Reduce::*;
import TLM3Stream::*;
import TLM3Utils::*;
import BusSwitch::*;


////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export TLM3Api::*;
export TLM3BRAM::*;
export TLM3CBusAdapter::*;
export TLM3Defines::*;
export TLM3Limit::*;
export TLM3Reorder::*;
export TLM3FlowControl::*;
export TLM3Ram::*;
export TLM3ReadWriteRam::*;
export TLM3Reduce::*;
export TLM3Stream::*;
export TLM3Utils::*;
export BusSwitch::*;

endpackage
