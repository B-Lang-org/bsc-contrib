package GenCRepr where

import List

type ByteList = List (Bit 8)

class ConvByteList n where
  toByteList :: Bit n -> ByteList
  fromByteList :: ByteList -> Bit n

instance ConvByteList 0 where
  toByteList _ = Nil
  fromByteList _ = 0

instance (Add 8 m n, ConvByteList m) => ConvByteList n where
  toByteList bs =
    case split bs of
      (h, t) -> h :> toByteList t
  fromByteList (Cons h t) = h ++ fromByteList t
  fromByteList Nil = 0

numCBytes :: Integer -> Maybe Integer
numCBytes numBytes =
  if numBytes <= 1 then Just 1
  else if numBytes <= 2 then Just 2
  else if numBytes <= 4 then Just 4
  else if numBytes <= 8 then Just 8
  else Nothing

bitsToBytes :: Integer -> Integer
bitsToBytes b = (((b - 1) / 8) + 1)

genCIntType :: Bool -> Integer -> (String, String)
genCIntType signed numBytes =
  let prefix = if signed then "int" else "uint"
  in case numCBytes numBytes of
    Just b -> (prefix +++ integerToString (b * 8) +++ "_t", "")
    Nothing -> (prefix +++ "8_t", "[" +++ integerToString numBytes +++ "]")

genCIntPack :: Integer -> String -> String -> String
genCIntPack numBytes val buf =
  let shiftPack :: Integer -> String
      shiftPack n = if n >= numBytes then "" else
           "**" +++ buf +++ " = 0xFF & (" +++ val +++ " >> " +++ integerToString (8 * (numBytes - n - 1)) +++ "); (*" +++ buf +++ ")++; " +++ shiftPack (n + 1)
  in case numCBytes numBytes of
    Just _ -> shiftPack 0
    Nothing ->
      "memcpy(*" +++ buf +++ ", &" +++ val +++ ", " +++ integerToString numBytes +++ "); " +++
      "*" +++ buf +++ " += " +++ integerToString numBytes +++ ";"

genCIntUnpack :: Integer -> String -> String -> String
genCIntUnpack numBytes val buf =
  let shiftUnpack :: Integer -> String
      shiftUnpack n =
        "((*" +++ buf +++ ")[" +++ integerToString n +++ "] << " +++ integerToString (8 * (numBytes - n - 1)) +++ ")" +++
        if n >= numBytes - 1 then "" else " | " +++ shiftUnpack (n + 1)
  in (case numCBytes numBytes of
        Just _ -> val +++ " = " +++ shiftUnpack 0 +++ ";"
        Nothing -> "memcpy(&" +++ val +++ ", *" +++ buf +++ ", " +++ integerToString numBytes +++ "); "
     ) +++ " *" +++ buf +++ " += " +++ integerToString numBytes +++ ";"

class GenCRepr a n | a -> n where
  genCType :: a -> (String, String)

  genCTypeDecl :: a -> Maybe String
  genCTypeDecl _ = Nothing

  pack :: a -> ByteList

  genCPack :: a -> String -> String -> String

  genCPackDecl :: a -> Maybe (String, String)
  genCPackDecl _ = Nothing

  unpack :: ByteList -> (a, ByteList)

  genCUnpack :: a -> String -> String -> String

  genCUnpackDecl :: a -> Maybe (String, String)
  genCUnpackDecl _ = Nothing

instance (ConvByteList b, Div b 8 n) => GenCRepr (UInt b) n where
  genCType _ = genCIntType False (valueOf n)

  pack x = toByteList $ Prelude.pack x
  genCPack _ = genCIntPack (valueOf n)

  unpack x = (Prelude.unpack $ fromByteList $ take (valueOf n) x, drop (valueOf n) x)
  genCUnpack _ = genCIntUnpack (valueOf n)

instance (ConvByteList b, Div b 8 n) => GenCRepr (Int b) n where
  genCType _ = genCIntType True (valueOf n)

  pack x = toByteList $ Prelude.pack x
  genCPack _ = genCIntPack (valueOf n)

  unpack x = (Prelude.unpack $ fromByteList $ take (valueOf n) x, drop (valueOf n) x)
  genCUnpack _ = genCIntUnpack (valueOf n)

instance GenCRepr Bool 1 where
  genCType _ = ("_Bool", "")

  pack x = zeroExtend (Prelude.pack x) :> Nil
  genCPack _ = genCIntPack 1

  unpack x = (Prelude.unpack $ truncate $ head x, tail x)
  genCUnpack _ = genCIntUnpack 1

instance (Generic a r, GenCRepr' r n) => GenCRepr a n where
  genCType _ = genCType' (_ :: r)
  genCTypeDecl _ = genCTypeDecl' (_ :: r)

  pack x = pack' $ from x
  genCPack _ = genCPack' (_ :: r)
  genCPackDecl _ = genCPackDecl' (_ :: r)

  unpack x =
    case unpack' x of
      (res, extra) -> (to res, extra)
  genCUnpack _ = genCUnpack' (_ :: r)
  genCUnpackDecl _ = genCUnpackDecl' (_ :: r)

class GenCRepr' a n | a -> n where
  genCType' :: a -> (String, String)
  genCTypeDecl' :: a -> Maybe String

  pack' :: a -> ByteList
  genCPack' :: a -> String -> String -> String
  genCPackDecl' :: a -> Maybe (String, String)

  unpack' :: ByteList -> (a, ByteList)
  genCUnpack' :: a -> String -> String -> String
  genCUnpackDecl' :: a -> Maybe (String, String)

-- Represent primitives as unsigned integers by default
instance (Bits a numBits, Div numBits 8 n, Mul n 8 numBitsPadded,
          Add numBits numPad numBitsPadded, ConvByteList numBitsPadded) =>
         GenCRepr' (ConcPrim a) n where
  genCType' _ = genCIntType False (valueOf n)
  genCTypeDecl' _ = Nothing

  pack' (ConcPrim x) = toByteList $ ((Prelude.pack x ++ 0) :: Bit numBitsPadded)
  genCPack' _ = genCIntPack (valueOf n)
  genCPackDecl' _ = Nothing

  unpack' x =
    (ConcPrim $ Prelude.unpack (split ((fromByteList $ take (valueOf n) x) :: Bit numBitsPadded)).fst,
     drop (valueOf n) x)
  genCUnpack' _ = genCIntUnpack (valueOf n)
  genCUnpackDecl' _ = Nothing

instance (GenCStructBody bodyRepr n) =>
         GenCRepr' (Meta (MetaData name pkg 1) (Meta (MetaConsNamed cName cIdx numFields) bodyRepr)) n where
  genCType' _ = (stringOf name, "")
  genCTypeDecl' _ = Just $ "typedef struct " +++ stringOf name +++ " {\n" +++
    genCStructBody (_ :: bodyRepr) False +++
    "} " +++ stringOf name +++ ";"

  pack' (Meta (Meta y)) = packStructBody y

  genCPack' _ val buf = "pack_" +++ stringOf name +++ "(" +++ val +++ ", " +++ buf +++ ");"

  genCPackDecl' _ = Just (
    "void pack_" +++ stringOf name +++ "(" +++ stringOf name +++ " val, uint8_t **buf);",
    "void pack_" +++ stringOf name +++ "(" +++ stringOf name +++ " val, uint8_t **buf) {\n" +++
    genCPackStructBody (_ :: bodyRepr) False "" +++
    "}")

  unpack' x =
    case unpackStructBody x of
      (res, extra) -> (Meta $ Meta res, extra)

  genCUnpack' _ val buf = val +++ " = unpack_" +++ stringOf name +++ "(" +++ buf +++ ");"

  genCUnpackDecl' _ = Just (
    stringOf name +++ " unpack_" +++ stringOf name +++ "(uint8_t **buf);",
    stringOf name +++ " unpack_" +++ stringOf name +++ "(uint8_t **buf) {\n" +++
    "\t" +++ stringOf name +++ " val;\n" +++
    genCUnpackStructBody (_ :: bodyRepr) False "" +++
    "\treturn val;\n" +++
    "}")

instance (GenCUnionBody tagBytes bodyRepr 0 bodyBytes,
          Log numCtors tagBits, Div tagBits 8 tagBytes, Add tagBytes bodyBytes n) =>
         GenCRepr' (Meta (MetaData name pkg numCtors) bodyRepr) n where
  genCType' _ = (stringOf name, "")
  genCTypeDecl' _ = Just $ "typedef struct " +++ stringOf name +++ " {\n" +++
    "\tenum " +++ stringOf name +++ "_tag { " +++
    genCEnumBody (_ :: Bit tagBytes) (_ :: bodyRepr) (stringOf name) +++
    " } tag;\n" +++
    "\tunion " +++ stringOf name +++ "_contents {\n" +++
    genCUnionBody (_ :: Bit tagBytes) (_ :: bodyRepr) (stringOf name) +++
    "\t} contents;\n" +++
    "} " +++ stringOf name +++ ";"

  pack' (Meta y) = packUnionBody (_ :: Bit tagBytes) y

  genCPack' _ val buf = "pack_" +++ stringOf name +++ "(" +++ val +++ ", " +++ buf +++ ");"

  genCPackDecl' _ = Just (
    "void pack_" +++ stringOf name +++ "(" +++ stringOf name +++ " val, uint8_t **buf);",
    "void pack_" +++ stringOf name +++ "(" +++ stringOf name +++ " val, uint8_t **buf) {\n" +++
    "\t" +++ genCIntPack (valueOf tagBytes) "val.tag" "buf" +++ "\n" +++
    "\t" +++ genCPackUnionBody (_ :: Bit tagBytes) (_ :: bodyRepr) (stringOf name) +++ " // Invalid tag, do nothing\n" +++
    "}")

  unpack' x =
    case unpackUnionBody (_ :: Bit tagBytes) x of
      (res, extra) -> (Meta res, extra)

  genCUnpack' _ val buf = val +++ " = unpack_" +++ stringOf name +++ "(" +++ buf +++ ");"

  genCUnpackDecl' _ = Just (
    stringOf name +++ " unpack_" +++ stringOf name +++ "(uint8_t **buf);",
    stringOf name +++ " unpack_" +++ stringOf name +++ "(uint8_t **buf) {\n" +++
    "\t" +++ stringOf name +++ " val;\n" +++
    "\t" +++ genCIntUnpack (valueOf tagBytes) "val.tag" "buf" +++ "\n" +++
    "\t" +++ genCUnpackUnionBody (_ :: Bit tagBytes) (_ :: bodyRepr) (stringOf name) +++ " // Invalid tag, do nothing\n" +++
    "\treturn val;\n" +++
    "}")

class GenCUnionBody nt a i n | nt a -> i n where
  genCEnumBody :: Bit nt -> a -> String -> String
  genCUnionBody :: Bit nt -> a -> String -> String

  packUnionBody :: Bit nt -> a -> ByteList
  genCPackUnionBody :: Bit nt -> a -> String -> String

  unpackUnionBody :: Bit nt -> ByteList -> (a, ByteList)
  genCUnpackUnionBody :: Bit nt -> a -> String -> String

instance (GenCUnionBody tagBytes a i1 n1, GenCUnionBody tagBytes b i2 n2,
          Max n1 n2 n,
          Mul tagBytes 8 tagBits, ConvByteList tagBits) =>
         GenCUnionBody tagBytes (Either a b) i1 n where
  genCEnumBody _ _ typeName =
    genCEnumBody (_ :: Bit tagBytes) (_ :: a) typeName +++ ", " +++
    genCEnumBody (_ :: Bit tagBytes) (_ :: b) typeName
  genCUnionBody _ _ typeName =
    genCUnionBody (_ :: Bit tagBytes) (_ :: a) typeName +++
    genCUnionBody (_ :: Bit tagBytes) (_ :: b) typeName

  packUnionBody _ (Left x) = packUnionBody (_ :: Bit tagBytes) x
  packUnionBody _ (Right x) = packUnionBody (_ :: Bit tagBytes) x
  genCPackUnionBody _ _ typeName =
    genCPackUnionBody (_ :: Bit tagBytes) (_ :: a) typeName +++ " else " +++
    genCPackUnionBody (_ :: Bit tagBytes) (_ :: b) typeName

  unpackUnionBody _ x =
    if fromByteList (take (valueOf tagBytes) x) == ((fromInteger (valueOf i1)) :: Bit tagBits)
    then case unpackUnionBody (_ :: Bit tagBytes) x of
      (res, extra) -> (Left res, extra)
    else case unpackUnionBody (_ :: Bit tagBytes) x of
      (res, extra) -> (Right res, extra)
  genCUnpackUnionBody _ _ typeName =
    genCUnpackUnionBody (_ :: Bit tagBytes) (_ :: a) typeName +++ " else " +++
    genCUnpackUnionBody (_ :: Bit tagBytes) (_ :: b) typeName

instance (GenCStructBody bodyRepr bodyBytes,
          Add tagBytes bodyBytes n, Mul tagBytes 8 tagBits, ConvByteList tagBits) =>
         GenCUnionBody tagBytes (Meta (MetaConsNamed ctorName ctorIdx numFields) bodyRepr) ctorIdx n where
  genCEnumBody _ _ typeName = typeName +++ "_" +++ stringOf ctorName
  genCUnionBody _ _ typeName =
    "\t\tstruct " +++ typeName +++ "_" +++ stringOf ctorName +++ " {\n" +++
    genCStructBody (_ :: bodyRepr) True +++
    "\t\t} " +++ stringOf ctorName +++ ";\n"

  packUnionBody _ (Meta x) =
    append (toByteList (Prelude.pack ((fromInteger $ valueOf ctorIdx) :: UInt tagBits))) $ packStructBody x
  genCPackUnionBody _ _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    genCPackStructBody (_ :: bodyRepr) True (".contents." +++ stringOf ctorName) +++ "\n" +++
    "\t}"

  unpackUnionBody _ x =
    case unpackStructBody $ drop (valueOf tagBytes) x of
      (res, extra) -> (Meta res, extra)
  genCUnpackUnionBody _ _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    genCUnpackStructBody (_ :: bodyRepr) True (".contents." +++ stringOf ctorName) +++ "\n" +++
    "\t}"

instance (GenCStructBody bodyRepr bodyBytes,
          Add tagBytes bodyBytes n, Mul tagBytes 8 tagBits, ConvByteList tagBits) =>
         GenCUnionBody tagBytes (Meta (MetaConsAnon ctorName ctorIdx numFields) bodyRepr) ctorIdx n where
  genCEnumBody _ _ typeName = typeName +++ "_" +++ stringOf ctorName
  genCUnionBody _ _ typeName =
    "\t\tstruct " +++ typeName +++ "_" +++ stringOf ctorName +++ " {\n" +++
    genCStructBody (_ :: bodyRepr) True +++
    "\t\t} " +++ stringOf ctorName +++ ";\n"

  packUnionBody _ (Meta x) =
    append (toByteList (Prelude.pack ((fromInteger $ valueOf ctorIdx) :: UInt tagBits))) $ packStructBody x
  genCPackUnionBody _ _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    genCPackStructBody (_ :: bodyRepr) True (".contents." +++ stringOf ctorName) +++ "\n" +++
    "\t}"

  unpackUnionBody _ x =
    case unpackStructBody $ drop (valueOf tagBytes) x of
      (res, extra) -> (Meta res, extra)
  genCUnpackUnionBody _ _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    genCUnpackStructBody (_ :: bodyRepr) True (".contents." +++ stringOf ctorName) +++ "\n" +++
    "\t}"

instance (GenCRepr a fieldBytes, Add tagBytes fieldBytes n, Mul tagBytes 8 tagBits, ConvByteList tagBits) =>
         GenCUnionBody tagBytes (Meta (MetaConsAnon ctorName ctorIdx 1) (Meta (MetaField fieldName fieldIdx) (Conc a))) ctorIdx n where
  genCEnumBody _ _ typeName = typeName +++ "_" +++ stringOf ctorName
  genCUnionBody _ _ _ =
    let (lType, rType) = genCType (_ :: a)
    in "\t\t" +++ lType +++ " " +++ stringOf ctorName +++ rType +++ ";\n"

  packUnionBody _ (Meta (Meta (Conc x))) =
    append (toByteList $ Prelude.pack ((fromInteger $ valueOf ctorIdx) :: UInt tagBits)) $ pack x
  genCPackUnionBody _ _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    "\t\t" +++ genCPack (_ :: a) ("val.contents." +++ stringOf ctorName) "buf" +++ "\n" +++
    "\t}"

  unpackUnionBody _ x =
    case unpack $ drop (valueOf tagBytes) x of
      (res, extra) -> (Meta $ Meta $ Conc res, extra)
  genCUnpackUnionBody _ _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    "\t\t" +++ genCUnpack (_ :: a) ("val.contents." +++ stringOf ctorName) "buf" +++ "\n" +++
    "\t}"


class GenCStructBody a n | a -> n where
  genCStructBody :: a -> Bool -> String
  packStructBody :: a -> ByteList
  genCPackStructBody :: a -> Bool -> String -> String
  unpackStructBody :: ByteList -> (a, ByteList)
  genCUnpackStructBody :: a -> Bool -> String -> String

instance (GenCStructBody a n1, GenCStructBody b n2,
          -- All data is byte-aligned for easier deserialization in C
          Div n1 8 n1Bytes, Mul n1Bytes 8 n1Padded, Add n1Padded n2 n,
          -- BSC isn't smart enough to infer this
          Add n1 n1Pad n1Padded) =>
         GenCStructBody (a, b) n where
  genCStructBody _ nested =
    genCStructBody (_ :: a) nested +++ genCStructBody (_ :: b) nested

  packStructBody (x, y) = packStructBody x `append` packStructBody y
  genCPackStructBody _ nested sel =
    genCPackStructBody (_ :: a) nested sel +++ genCPackStructBody (_ :: b) nested sel

  unpackStructBody x =
    case unpackStructBody x of
      (res1, extra1) ->
        case unpackStructBody extra1 of
          (res2, extra2) -> ((res1, res2), extra2)
  genCUnpackStructBody _ nested sel =
    genCUnpackStructBody (_ :: a) nested sel +++ genCUnpackStructBody (_ :: b) nested sel

instance GenCStructBody () 0 where
  genCStructBody _ _ = ""
  packStructBody () = Nil
  genCPackStructBody _ _ _ = ""
  unpackStructBody x = ((), x)
  genCUnpackStructBody _ _ _ = ""

instance (GenCRepr a n) => GenCStructBody (Meta (MetaField name idx) (Conc a)) n where
  genCStructBody _ nested =
    let (lType, rType) = genCType (_ :: a)
    in (if nested then "\t\t" else "") +++ "\t" +++ lType +++ " " +++ stringOf name +++ rType +++ ";\n"

  packStructBody (Meta (Conc x)) = pack x
  genCPackStructBody _ nested sel =
    (if nested then "\t" else "") +++
    "\t" +++ genCPack (_ :: a) ("val" +++ sel +++ "." +++ stringOf name) "buf" +++ "\n"

  unpackStructBody x =
    case unpack x of
      (res, extra) -> (Meta $ Conc res, extra)
  genCUnpackStructBody _ nested sel =
    (if nested then "\t" else "") +++
    "\t" +++ genCUnpack (_ :: a) ("val" +++ sel +++ "." +++ stringOf name) "buf" +++ "\n"


-- Helper to allow a tuple of types to be all easily translated together
class GenCDecls a where
  genCHeaderDecls :: a -> String
  genCImplDecls :: a -> String

instance (GenCDecls a, GenCDecls b) => GenCDecls (a, b) where
  genCHeaderDecls _ = genCHeaderDecls (_ :: a) +++ genCHeaderDecls (_ :: b)
  genCImplDecls _ = genCImplDecls (_ :: a) +++ genCImplDecls (_ :: b)

instance GenCDecls () where
  genCHeaderDecls _ = ""
  genCImplDecls _ = ""

instance (GenCRepr a n) => GenCDecls a where
  genCHeaderDecls p =
    (case genCTypeDecl p of
        Just d -> d +++ "\n"
        Nothing -> ""
    ) +++
    (case genCPackDecl p of
       Just (d, _) -> d +++ "\n"
       Nothing -> ""
    ) +++
    (case genCUnpackDecl p of
       Just (d, _) -> d +++ "\n\n"
       Nothing -> ""
    )

  genCImplDecls p =
    (case genCPackDecl p of
       Just (_, d) -> d +++ "\n\n"
       Nothing -> ""
    ) +++
    (case genCUnpackDecl p of
       Just (_, d) -> d +++ "\n\n"
       Nothing -> ""
    )

-- Driver to all write C declarations for some types
writeCDecls :: (GenCDecls tys) => String -> tys -> Module Empty
writeCDecls baseName proxy = do
  let headerName = (baseName +++ ".h")
  let implName = (baseName +++ ".c")
  let headerContents =
        "#include <stdint.h>\n\n\n" +++
        genCHeaderDecls proxy
  let implContents =
        "#include <stdlib.h>\n#include <string.h>\n\n#include \"" +++ headerName +++ "\"\n\n\n" +++
        genCImplDecls proxy
  stdout <- openFile "/dev/stdout" WriteMode
  h <- openFile headerName WriteMode
  hPutStr h headerContents
  hClose h
  hPutStrLn stdout ("Header file created: " +++ headerName)
  c <- openFile implName WriteMode
  hPutStr c implContents
  hClose c
  hPutStrLn stdout ("C implementation file created: " +++ implName)
  hClose stdout
