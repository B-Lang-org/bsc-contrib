// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause

package Axi;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AxiDefines::*;
import AxiExtend::*;
import AxiMaster::*;
import AxiSlave::*;
import AxiRdBus::*;
import AxiWrBus::*;
import AxiPC::*;
// import AxiMonitor::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AxiDefines::*;
export AxiExtend::*;
export AxiMaster::*;
export AxiSlave::*;
export AxiRdBus::*;
export AxiWrBus::*;
export AxiPC::*;
// export AxiMonitor::*;

endpackage
