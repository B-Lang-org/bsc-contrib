
import "BDPI" function ActionValue#(Bit#(48)) getInstr();
import "BDPI" function Action putResult(Bit#(48) res);

