// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause

package Axi4;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import Axi4Defines::*;
import Axi4Master::*;
import Axi4Slave::*;
import Axi4PC::*;

import Axi4LDefines::*;
import Axi4LMaster::*;
import Axi4LSlave::*;
import Axi4LPC::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export Axi4Defines::*;
export Axi4Master::*;
export Axi4Slave::*;
export Axi4PC::*;

export Axi4LDefines::*;
export Axi4LMaster::*;
export Axi4LSlave::*;
export Axi4LPC::*;

endpackage
