// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause

package DDR2;

import DDR2Types::*;
import DDR2FakeBurst::*;
import ML507_DDR2::*;
import ML507_mig_33_wrapper::*;

export DDR2Types::*;
export DDR2FakeBurst::*;
export ML507_DDR2::*;
export ML507_mig_33_wrapper::*;

endpackage
