////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause
//
////////////////////////////////////////////////////////////////////////////////
//  Filename      : Xilinx.bsv
//  Description   : Xilinx specific libraries
////////////////////////////////////////////////////////////////////////////////
package Xilinx;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import XilinxCells       ::*;
import XilinxClocks      ::*;
import XilinxUtils       ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export XilinxCells       ::*;
import XilinxClocks      ::*;
export XilinxUtils       ::*;

endpackage: Xilinx
