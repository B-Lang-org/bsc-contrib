package GenCRepr where

numCBytes :: Integer -> Maybe Integer
numCBytes numBits =
  if numBits <= 8 then Just 1
  else if numBits <= 16 then Just 2
  else if numBits <= 32 then Just 4
  else if numBits <= 64 then Just 8
  else Nothing

bitsToBytes :: Integer -> Integer
bitsToBytes b = (((b - 1) / 8) + 1)

genCIntType :: Bool -> Integer -> (String, String)
genCIntType signed numBits =
  let prefix = if signed then "int" else "uint"
  in case numCBytes numBits of
    Just b -> (prefix +++ integerToString (b * 8) +++ "_t", "")
    Nothing -> (prefix +++ "8_t", "[" +++ integerToString (bitsToBytes numBits) +++ "]")

genCIntPack :: Integer -> String -> String -> String
genCIntPack numBits val buf =
  let numBytes = bitsToBytes numBits
      shiftPack :: Integer -> String
      shiftPack n = if n >= numBytes then "" else
           "**" +++ buf +++ " = 0xFF & (" +++ val +++ " >> " +++ integerToString (8 * (numBytes - n - 1)) +++ "); (*" +++ buf +++ ")++; " +++ shiftPack (n + 1)
  in case numCBytes numBits of
    Just _ -> shiftPack 0
    Nothing ->
      "memcpy(*" +++ buf +++ ", &" +++ val +++ ", " +++ integerToString numBytes +++ "); " +++
      "*" +++ buf +++ " += " +++ integerToString numBytes +++ ";"

genCIntUnpack :: Integer -> String -> String -> String
genCIntUnpack numBits val buf =
  let numBytes = bitsToBytes numBits
      shiftUnpack :: Integer -> String
      shiftUnpack n =
        "((*" +++ buf +++ ")[" +++ integerToString n +++ "] << " +++ integerToString (8 * (numBytes - n - 1)) +++ ")" +++
        if n >= numBytes - 1 then "" else " | " +++ shiftUnpack (n + 1)
  in (case numCBytes numBits of
        Just _ -> val +++ " = " +++ shiftUnpack 0 +++ ";"
        Nothing -> "memcpy(&" +++ val +++ ", *" +++ buf +++ ", " +++ integerToString numBytes +++ "); "
     ) +++ " *" +++ buf +++ " += " +++ integerToString numBytes +++ ";"

class GenCRepr a n | a -> n where
  genCType :: a -> (String, String)

  genCTypeDecl :: a -> Maybe String
  genCTypeDecl _ = Nothing

  pack :: a -> Bit n

  genCPack :: a -> String -> String -> String

  genCPackDecl :: a -> Maybe (String, String)
  genCPackDecl _ = Nothing

  unpack :: Bit n -> a

  genCUnpack :: a -> String -> String -> String

  genCUnpackDecl :: a -> Maybe (String, String)
  genCUnpackDecl _ = Nothing

instance GenCRepr (UInt n) n where
  genCType _ = genCIntType False (valueOf n)

  pack = Prelude.pack
  genCPack _ = genCIntPack (valueOf n)

  unpack = Prelude.unpack
  genCUnpack _ = genCIntUnpack (valueOf n)

instance GenCRepr (Int n) n where
  genCType _ = genCIntType True (valueOf n)

  pack = Prelude.pack
  genCPack _ = genCIntPack (valueOf n)

  unpack = Prelude.unpack
  genCUnpack _ = genCIntUnpack (valueOf n)

-- Booleans are each packed as an entire byte, for now
instance GenCRepr Bool 8 where
  genCType _ = ("_Bool", "")

  pack x = extend $ Prelude.pack x
  genCPack _ = genCIntPack 1

  unpack x = Prelude.unpack $ truncate x
  genCUnpack _ = genCIntUnpack 1

instance (Generic a r, GenCRepr' a r n) => GenCRepr a n where
  genCType p = genCType' p ((from p) :: r)
  genCTypeDecl p = genCTypeDecl' p ((from p) :: r)
  pack = pack' ((error "proxy") :: r)
  genCPack p = genCPack' p ((from p) :: r)
  genCPackDecl p = genCPackDecl' p ((from p) :: r)
  unpack = unpack' ((error "proxy") :: r)
  genCUnpack p = genCUnpack' p ((from p) :: r)
  genCUnpackDecl p = genCUnpackDecl' p ((from p) :: r)

-- Helper type class for coherent dispach on generic representation
class GenCRepr' a r n | a r -> n where
  genCType' :: a -> r -> (String, String)
  genCTypeDecl' :: a -> r -> Maybe String

  pack' :: r -> a -> Bit n
  genCPack' :: a -> r -> String -> String -> String
  genCPackDecl' :: a -> r -> Maybe (String, String)

  unpack' :: r -> Bit n -> a
  genCUnpack' :: a -> r -> String -> String -> String
  genCUnpackDecl' :: a -> r -> Maybe (String, String)

-- Default: serialize to Bits representation and pack as an integer
instance (Generic a r, Bits a n) => GenCRepr' a r n where
  genCType' _ _ = genCIntType False (valueOf n)
  genCTypeDecl' _ _ = Nothing

  pack' _ = Prelude.pack
  genCPack' _ _ = genCIntPack (valueOf n)
  genCPackDecl' _ _ = Nothing

  unpack' _ = Prelude.unpack
  genCUnpack' _ _ = genCIntUnpack (valueOf n)
  genCUnpackDecl' _ _ = Nothing

instance (Generic a (Meta (MetaData name pkg 1) (Meta (MetaConsNamed cName cIdx numFields) bodyRepr)),
          GenCStructBody bodyRepr n) =>
         GenCRepr' a (Meta (MetaData name pkg 1) (Meta (MetaConsNamed cName cIdx numFields) bodyRepr)) n where
  genCType' _ _ = (stringOf name, "")
  genCTypeDecl' _ _ = Just $ "typedef struct " +++ stringOf name +++ " {\n" +++
    genCStructBody ((error "proxy") :: bodyRepr) False +++
    "} " +++ stringOf name +++ ";"

  pack' _ x =
    case from x of
      (Meta (Meta y)) -> packStructBody y

  genCPack' _ _ val buf = "pack_" +++ stringOf name +++ "(" +++ val +++ ", " +++ buf +++ ");"

  genCPackDecl' _ _ = Just (
    "void pack_" +++ stringOf name +++ "(" +++ stringOf name +++ " val, uint8_t **buf);",
    "void pack_" +++ stringOf name +++ "(" +++ stringOf name +++ " val, uint8_t **buf) {\n" +++
    genCPackStructBody ((error "proxy") :: bodyRepr) False "" +++
    "}")

  unpack' _ x = to $ Meta $ Meta $ unpackStructBody x

  genCUnpack' _ _ val buf = val +++ " = unpack_" +++ stringOf name +++ "(" +++ buf +++ ");"

  genCUnpackDecl' _ _ = Just (
    stringOf name +++ " unpack_" +++ stringOf name +++ "(uint8_t **buf);",
    stringOf name +++ " unpack_" +++ stringOf name +++ "(uint8_t **buf) {\n" +++
    "\t" +++ stringOf name +++ " val;\n" +++
    genCUnpackStructBody ((error "proxy") :: bodyRepr) False "" +++
    "\treturn val;\n" +++
    "}")

instance (Generic a (Meta (MetaData name pkg numCtors) bodyRepr),
          GenCUnionBody 0 bodyRepr n,
          -- For simplicity the tag must fit in a single byte, for now.
          Add 8 bodyBits n, Max numCtors 255 255) =>
         GenCRepr' a (Meta (MetaData name pkg numCtors) bodyRepr) n where
  genCType' _ _ = (stringOf name, "")
  genCTypeDecl' _ _ = Just $ "typedef struct " +++ stringOf name +++ " {\n" +++
    "\tenum " +++ stringOf name +++ "_tag { " +++
    genCEnumBody ((error "proxy") :: bodyRepr) (stringOf name) +++
    " } tag;\n" +++
    "\tunion " +++ stringOf name +++ "_contents {\n" +++
    genCUnionBody ((error "proxy") :: bodyRepr) (stringOf name) +++
    "\t} contents;\n" +++
    "} " +++ stringOf name +++ ";"

  pack' _ x =
    case from x of
      (Meta y) -> packUnionBody y

  genCPack' _ _ val buf = "pack_" +++ stringOf name +++ "(" +++ val +++ ", " +++ buf +++ ");"

  genCPackDecl' _ _ = Just (
    "void pack_" +++ stringOf name +++ "(" +++ stringOf name +++ " val, uint8_t **buf);",
    "void pack_" +++ stringOf name +++ "(" +++ stringOf name +++ " val, uint8_t **buf) {\n" +++
    "\t**buf = val.tag; (*buf)++;\n" +++
    "\t" +++ genCPackUnionBody ((error "proxy") :: bodyRepr) (stringOf name) +++ " // Invalid tag, do nothing\n" +++
    "}")

  unpack' _ x = to $ Meta $ uncurry unpackUnionBody $ split x

  genCUnpack' _ _ val buf = val +++ " = unpack_" +++ stringOf name +++ "(" +++ buf +++ ");"

  genCUnpackDecl' _ _ = Just (
    stringOf name +++ " unpack_" +++ stringOf name +++ "(uint8_t **buf);",
    stringOf name +++ " unpack_" +++ stringOf name +++ "(uint8_t **buf) {\n" +++
    "\t" +++ stringOf name +++ " val;\n" +++
    "\tval.tag = **buf; (*buf)++;\n" +++
    "\t" +++ genCUnpackUnionBody ((error "proxy") :: bodyRepr) (stringOf name) +++ " // Invalid tag, do nothing\n" +++
    "\treturn val;\n" +++
    "}")

class GenCUnionBody i a n | a -> i n where
  genCEnumBody :: a -> String -> String
  genCUnionBody :: a -> String -> String

  packUnionBody :: a -> Bit n
  genCPackUnionBody :: a -> String -> String

  unpackUnionBody :: (Add 8 m n) => Bit 8 -> Bit m -> a
  genCUnpackUnionBody :: a -> String -> String

instance (Add i 1 i2,
          GenCUnionBody i a n1, GenCUnionBody i2 b n2,
          Max n1 n2 n,
          Add 8 m1 n1, Add 8 m2 n2, Add m1 m1Pad n, Add m2 m2Pad n,
          Add n1 n1Pad n, Add n2 n2Pad n) =>
         GenCUnionBody i (Either a b) n where
  genCEnumBody _ typeName =
    genCEnumBody ((error "proxy") :: a) typeName +++ ", " +++ genCEnumBody ((error "proxy") :: b) typeName
  genCUnionBody _ typeName =
    genCUnionBody ((error "proxy") :: a) typeName +++ genCUnionBody  ((error "proxy") :: b) typeName

  packUnionBody (Left x) = packUnionBody x ++ fromInteger 0
  packUnionBody (Right x) = packUnionBody x ++ fromInteger 0
  genCPackUnionBody _ typeName =
    genCPackUnionBody ((error "proxy") :: a) typeName +++ " else " +++ genCPackUnionBody  ((error "proxy") :: b) typeName

  unpackUnionBody tag body =
    if tag == fromInteger (valueOf i)
    then Left $ unpackUnionBody tag ((split body).fst :: Bit n1)
    else Right $ unpackUnionBody tag ((split body).fst :: Bit n2)
  genCUnpackUnionBody _ typeName =
    genCUnpackUnionBody ((error "proxy") :: a) typeName +++ " else " +++ genCUnpackUnionBody  ((error "proxy") :: b) typeName

instance (GenCStructBody bodyRepr bodyBits, Add 8 bodyBits n) =>
         GenCUnionBody i (Meta (MetaConsNamed ctorName ctorIdx numFields) bodyRepr) n where
  genCEnumBody _ typeName = typeName +++ "_" +++ stringOf ctorName
  genCUnionBody _ typeName =
    "\t\tstruct " +++ typeName +++ "_" +++ stringOf ctorName +++ " {\n" +++
    genCStructBody ((error "proxy") :: bodyRepr) True +++
    "\t\t} " +++ stringOf ctorName +++ ";\n"

  packUnionBody (Meta x) = Prelude.pack ((fromInteger $ valueOf ctorIdx) :: UInt 8) ++ packStructBody x
  genCPackUnionBody _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    genCPackStructBody ((error "proxy") :: bodyRepr) True (".contents." +++ stringOf ctorName) +++ "\n" +++
    "\t}"

  genCUnpackUnionBody _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    genCUnpackStructBody ((error "proxy") :: bodyRepr) True (".contents." +++ stringOf ctorName) +++ "\n" +++
    "\t}"

instance (GenCStructBody bodyRepr bodyBits, Add 8 bodyBits n) =>
         GenCUnionBody i (Meta (MetaConsAnon ctorName ctorIdx numFields) bodyRepr) n where
  genCEnumBody _ typeName = typeName +++ "_" +++ stringOf ctorName
  genCUnionBody _ typeName =
    "\t\tstruct " +++ typeName +++ "_" +++ stringOf ctorName +++ " {\n" +++
    genCStructBody ((error "proxy") :: bodyRepr) True +++
    "\t\t} " +++ stringOf ctorName +++ ";\n"

  packUnionBody (Meta x) = Prelude.pack ((fromInteger $ valueOf ctorIdx) :: UInt 8) ++ packStructBody x
  genCPackUnionBody _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    genCPackStructBody ((error "proxy") :: bodyRepr) True (".contents." +++ stringOf ctorName) +++ "\n" +++
    "\t}"

  genCUnpackUnionBody _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    genCUnpackStructBody ((error "proxy") :: bodyRepr) True (".contents." +++ stringOf ctorName) +++ "\n" +++
    "\t}"

instance (GenCRepr a fieldBits, Add 8 fieldBits n) =>
         GenCUnionBody i (Meta (MetaConsAnon ctorName ctorIdx 1) (Meta (MetaField fieldName fieldIdx) (Conc a))) n where
  genCEnumBody _ typeName = typeName +++ "_" +++ stringOf ctorName
  genCUnionBody _ _ =
    let (lType, rType) = genCType ((error "proxy") :: a)
    in "\t\t" +++ lType +++ " " +++ stringOf ctorName +++ rType +++ ";\n"

  packUnionBody (Meta (Meta (Conc x))) = Prelude.pack ((fromInteger $ valueOf ctorIdx) :: UInt 8) ++ pack x
  genCPackUnionBody _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    "\t\t" +++ genCPack ((error "proxy") :: a) ("val.contents." +++ stringOf ctorName) "buf" +++ "\n" +++
    "\t}"

  genCUnpackUnionBody _ typeName =
    "if (val.tag == " +++ typeName +++ "_" +++ stringOf ctorName +++ ") {\n" +++
    "\t\t" +++ genCUnpack ((error "proxy") :: a) ("val.contents." +++ stringOf ctorName) "buf" +++ "\n" +++
    "\t}"


class GenCStructBody a n | a -> n where
  genCStructBody :: a -> Bool -> String
  packStructBody :: a -> Bit n
  genCPackStructBody :: a -> Bool -> String -> String
  unpackStructBody :: Bit n -> a
  genCUnpackStructBody :: a -> Bool -> String -> String

instance (GenCStructBody a n1, GenCStructBody b n2,
          -- All data is byte-aligned for easier deserialization in C
          Div n1 8 n1Bytes, Mul n1Bytes 8 n1Padded, Add n1Padded n2 n,
          -- BSC isn't smart enough to infer this
          Add n1 n1Pad n1Padded) =>
         GenCStructBody (a, b) n where
  genCStructBody _ nested =
    genCStructBody ((error "proxy") :: a) nested +++ genCStructBody ((error "proxy") :: b) nested

  packStructBody (x, y) = zeroExtend (packStructBody x) ++ packStructBody y
  genCPackStructBody _ nested sel =
    genCPackStructBody ((error "proxy") :: a) nested sel +++ genCPackStructBody ((error "proxy") :: b) nested sel

  unpackStructBody bs =
    let (xbs, ybs) = (split bs) :: (Bit n1Padded, Bit n2)
    in (unpackStructBody $ truncate xbs, unpackStructBody ybs)
  genCUnpackStructBody _ nested sel =
    genCUnpackStructBody ((error "proxy") :: a) nested sel +++ genCUnpackStructBody ((error "proxy") :: b) nested sel

instance GenCStructBody () 0 where
  genCStructBody _ _ = ""
  packStructBody () = 0'b0
  genCPackStructBody _ _ _ = ""
  unpackStructBody _ = ()
  genCUnpackStructBody _ _ _ = ""

instance (GenCRepr a n) => GenCStructBody (Meta (MetaField name idx) (Conc a)) n where
  genCStructBody _ nested =
    let (lType, rType) = genCType ((error "proxy") :: a)
    in (if nested then "\t\t" else "") +++ "\t" +++ lType +++ " " +++ stringOf name +++ rType +++ ";\n"

  packStructBody (Meta (Conc x)) = pack x
  genCPackStructBody _ nested sel =
    (if nested then "\t" else "") +++
    "\t" +++ genCPack ((error "proxy") :: a) ("val" +++ sel +++ "." +++ stringOf name) "buf" +++ "\n"

  unpackStructBody x = Meta $ Conc $ unpack x
  genCUnpackStructBody _ nested sel =
    (if nested then "\t" else "") +++
    "\t" +++ genCUnpack ((error "proxy") :: a) ("val" +++ sel +++ "." +++ stringOf name) "buf" +++ "\n"


-- Helper to allow a tuple of types to be all easily translated together
class GenCDecls a where
  genCHeaderDecls :: a -> String
  genCImplDecls :: a -> String

instance (GenCDecls a, GenCDecls b) => GenCDecls (a, b) where
  genCHeaderDecls _ = genCHeaderDecls ((error "proxy") :: a) +++ genCHeaderDecls ((error "proxy") :: b)
  genCImplDecls _ = genCImplDecls ((error "proxy") :: a) +++ genCImplDecls ((error "proxy") :: b)

instance GenCDecls () where
  genCHeaderDecls _ = ""
  genCImplDecls _ = ""

instance (GenCRepr a n) => GenCDecls a where
  genCHeaderDecls p =
    (case genCTypeDecl p of
        Just d -> d +++ "\n"
        Nothing -> ""
    ) +++
    (case genCPackDecl p of
       Just (d, _) -> d +++ "\n"
       Nothing -> ""
    ) +++
    (case genCUnpackDecl p of
       Just (d, _) -> d +++ "\n\n"
       Nothing -> ""
    )

  genCImplDecls p =
    (case genCPackDecl p of
       Just (_, d) -> d +++ "\n\n"
       Nothing -> ""
    ) +++
    (case genCUnpackDecl p of
       Just (_, d) -> d +++ "\n\n"
       Nothing -> ""
    )

-- Driver to all write C declarations for some types
writeCDecls :: (GenCDecls tys) => String -> tys -> Module Empty
writeCDecls baseName proxy = do
  let headerName = (baseName +++ ".h")
  let implName = (baseName +++ ".c")
  let headerContents =
        "#include <stdint.h>\n\n\n" +++
        genCHeaderDecls proxy
  let implContents =
        "#include <stdlib.h>\n#include <string.h>\n\n#include \"" +++ headerName +++ "\"\n\n\n" +++
        genCImplDecls proxy
  stdout <- openFile "/dev/stdout" WriteMode
  h <- openFile headerName WriteMode
  hPutStr h headerContents
  hClose h
  hPutStrLn stdout ("Header file created: " +++ headerName)
  c <- openFile implName WriteMode
  hPutStr c implContents
  hClose c
  hPutStrLn stdout ("C implementation file created: " +++ implName)
  hClose stdout
