
import "BDPI" function Bit#(32) test_fn(Bit#(48) arg);
     
