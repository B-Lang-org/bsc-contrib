package GenCRepr where

numCBytes :: Integer -> Maybe Integer
numCBytes numBits =
  if numBits < 8 then Just 1
  else if numBits < 16 then Just 2
  else if numBits < 32 then Just 4
  else if numBits < 64 then Just 8
  else Nothing

genCIntType :: Bool -> Integer -> (String, String)
genCIntType signed numBits =
  let prefix = if signed then "int" else "uint"
  in case numCBytes numBits of
    Just b -> (prefix +++ integerToString (b * 8) +++ "_t", "")
    Nothing -> (prefix +++ "8_t", "[" +++ integerToString (((numBits - 1) / 8) + 1) +++ "]")

class GenCRepr a where
  genCType :: a -> (String, String)
  
  genCTypeDecl :: a -> Maybe String
  genCTypeDecl _ = Nothing

  genCPack :: a -> Maybe (String, String)
  genCPack _ = Nothing

instance GenCRepr (Bit n) where
  genCType _ = genCIntType False (valueOf n)

instance GenCRepr (UInt n) where
  genCType _ = genCIntType False (valueOf n)

instance GenCRepr (Int n) where
  genCType _ = genCIntType True (valueOf n)

instance GenCRepr Bool where
  genCType _ = ("_Bool", "")

instance (Generic a (Meta (MetaData name pkg 1) (Meta (MetaConsNamed cName cIdx numFields) bodyRepr)),
          GenCStructBody bodyRepr) => GenCRepr a where
  genCType _ = (stringOf name, "")
  genCTypeDecl _ = Just $ "typedef struct " +++ stringOf name +++ " {\n" +++ genCStructBody ((error "proxy") :: bodyRepr) +++ "} " +++ stringOf name +++ ";"

class GenCStructBody a where
  genCStructBody :: a -> String

instance (GenCStructBody a, GenCStructBody b) => GenCStructBody (a, b) where
  genCStructBody _ = genCStructBody ((error "proxy") :: a) +++ genCStructBody ((error "proxy") :: b)

instance GenCStructBody () where
  genCStructBody _ = ""

instance (GenCRepr a) => GenCStructBody (Meta (MetaField name idx) (Conc a)) where
  genCStructBody _ =
    let (lType, rType) = genCType ((error "proxy") :: a)
    in "\t" +++ lType +++ " " +++ stringOf name +++ rType +++ ";\n"


-- Helper to allow a tuple of types to be all easily translated together
class GenCDecls a where
  genCTypeDecls :: a -> String

instance (GenCDecls a, GenCDecls b) => GenCDecls (a, b) where
  genCTypeDecls _ = genCTypeDecls ((error "proxy") :: a) +++ genCTypeDecls ((error "proxy") :: b)

instance GenCDecls () where
  genCTypeDecls _ = ""

instance (GenCRepr a) => GenCDecls a where
  genCTypeDecls p =
    case genCTypeDecl p of
      Just d -> d +++ "\n\n"
      Nothing -> ""

-- Driver to all write C declarations for some types
writeCDecls :: (GenCDecls tys) => String -> tys -> Module Empty
writeCDecls baseName proxy = do
  let typeDecls = genCTypeDecls proxy
  let headerName = (baseName +++ ".h")
  let implName = (baseName +++ ".c")
  let headerContents = "#include <stdint.h>\n\n\n" +++ typeDecls
  let implContents = "#include <stdlib.h>\n#include <string.h>\n\n#include \"" +++ headerName +++ "\"\n\n\n"
  stdout <- openFile "/dev/stdout" WriteMode
  h <- openFile headerName WriteMode
  hPutStr h headerContents
  hClose h
  hPutStrLn stdout ("Header file created: " +++ headerName)
  c <- openFile implName WriteMode
  hPutStr c implContents
  hClose c
  hPutStrLn stdout ("C implementation file created: " +++ implName)
  hClose stdout
