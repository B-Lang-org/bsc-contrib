// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause

package TLM;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import TLMCBusAdapter::*;
import TLMDefines::*;
import TLMRam::*;
import TLMReadWriteRam::*;
import TLMReduce::*;
import TLMUtils::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export TLMCBusAdapter::*;
export TLMDefines::*;
export TLMRam::*;
export TLMReadWriteRam::*;
export TLMReduce::*;
export TLMUtils::*;

endpackage
