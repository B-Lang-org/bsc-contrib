// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause

package AHB;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AHBArbiter::*;
import AHBBus::*;
import AHBDefines::*;
import AHBMaster::*;
import AHBPC::*;
import AHBSlave::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AHBArbiter::*;
export AHBBus::*;
export AHBDefines::*;
export AHBMaster::*;
export AHBPC::*;
export AHBSlave::*;

endpackage
