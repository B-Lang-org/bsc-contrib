
import "BDPI" function ActionValue#(Bool) messageAvailable();
import "BDPI" function ActionValue#(Bit#(56)) getMessage();
import "BDPI" function Action putMessage(Bit#(56) res);
