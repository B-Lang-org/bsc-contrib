package Counter where

import GenCRepr
import GenCMsg
import CounterIface
import CShow
import Vector

type Id = Bit 16 -- Try changing the size (will need to update in CounterIface.bsv)

-- Try adding/reordering constructors
data Command = Num { id :: Id; val :: Int 16; }
             | Reset (Int 16)
             | Halt
  deriving (Bits)

struct Result a =
  id :: Id
  val :: a
 deriving (Bits)

interface CounterMsgs =
  -- In order of highest to lowest urgency, try changing the order!
  commands :: Rx Command
  sums     :: Tx (Result (Int 16))
  products :: Tx (Result (Int 32))

{-# verilog mkCounter #-}
mkCounter :: Module Empty
mkCounter = module
  writeCMsgDecls "counter" (_ :: CounterMsgs)

  msgMgr <- mkMsgManager
  let msgs :: CounterMsgs = msgMgr.fifos

  sum :: Reg (Int 16) <- mkReg 0
  product :: Reg (Int 32) <- mkReg 1

  rules
    "handle_command": when True ==> do
      let c :: Command = msgs.commands.first
      msgs.commands.deq
      -- $display "Handling command " (cshow c)
      case c of
        Num { id = id; val = val; } -> do
          let newSum = sum + val
          let newProduct = product * signExtend val
          msgs.sums.enq (Result { id = id; val = newSum; })
          msgs.products.enq (Result { id = id; val = newProduct; })
          sum := newSum
          product := newProduct
        Reset val -> do
          sum := val
          product := signExtend val
        Halt -> $finish

    "recieve_message": when messageAvailable ==> do
      m <- getMessage
      let mBytes = unpack m
      -- $display "B recieved message " (cshow mBytes)
      msgMgr.putMsg mBytes

    "send_message": when True ==> do
      (_, mBytes) <- msgMgr.getMsg
      -- $display "B sending message " (cshow mBytes)
      putMessage (pack mBytes)
