// Copyright (c) 2020 Bluespec, Inc. All rights reserved.
//
// SPDX-License-Identifier: BSD-3-Clause

package Ahb;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AhbArbiter::*;
import AhbBus::*;
import AhbDefines::*;
import AhbMaster::*;
import AhbPC::*;
import AhbSlave::*;
import AhbToAhbBridge::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AhbArbiter::*;
export AhbBus::*;
export AhbDefines::*;
export AhbMaster::*;
export AhbPC::*;
export AhbSlave::*;
export AhbToAhbBridge::*;

endpackage
