
import "BDPI" function ActionValue#(Bit#(48)) test_fn(Bit#(64) arg);
     
